module logistic_regression (
    
);
    
endmodule