module matrix_memory (
    
);
    
endmodule