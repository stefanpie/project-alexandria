module support_vector_machine (
    
);
    
endmodule