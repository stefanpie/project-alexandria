module linear_regression (
    input data_i,
    input weights_i
);
    
endmodule