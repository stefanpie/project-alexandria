module decision_tree (
    
);
    
endmodule